// File: tb/common/pkg/common_pkg.sv
`ifndef COMMON_PKG_SV
`define COMMON_PKG_SV

package common_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"



endpackage: common_pkg

`endif // COMMON_PKG_SV
