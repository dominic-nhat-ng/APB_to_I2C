package apb_tests_pkg;
    import uvm_pkg::*;
    import apb_pkg::*;
    `include "uvm_macros.svh"
    `include "apb_tests/apb_base_test.sv"
endpackage
