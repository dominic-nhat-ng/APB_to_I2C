package i2c_tests_pkg;
    import uvm_pkg::*;
    import i2c_pkg::*;
    `include "uvm_macros.svh"
    `include "i2c_tests/i2c_base_test.sv"
endpackage
