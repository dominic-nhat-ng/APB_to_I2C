class apb_base_test extends uvm_test;

endclass
