package test_pkg;
    import uvm_pkg::*;
    import apb_pkg::*;
    import i2c_pkg::*;
    import apb_tests_pkg::*;
    import i2c_tests_pkg::*;
    `include "uvm_macros.svh"
endpackage
