`ifndef APB_PKG_SV
`define APB_PKG_SV

package apb_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "agent/apb_transaction.sv"
  `include "agent/apb_sequencer.sv"
  `include "agent/apb_driver.sv"
  `include "agent/apb_monitor.sv"
  `include "env/apb_agent.sv"
  `include "env/apb_scoreboard.sv"
  `include "env/apb_env.sv"
  `include "sequences/apb_base_sequence.sv"

endpackage: apb_pkg

`endif // APB_PKG_SV
